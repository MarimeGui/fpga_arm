package Utilities;

    bit [4:0] NOP = 5'd0;
    bit [4:0] ADD = 5'd1;
    bit [4:0] SUB = 5'd2;
    bit [4:0] AND = 5'd3;
    bit [4:0] EOR = 5'd4;
    bit [4:0] CMP = 5'd5;
    bit [4:0] LSL = 5'd6;
    bit [4:0] LSR = 5'd7;
    bit [4:0] MOV = 5'd8;
    bit [4:0] STR = 5'd9;
    bit [4:0] LDR = 5'd10;
    //bit [4:0] PUSH = 5'd11;
    //bit [4:0] POP = 5'd12;

    typedef struct packed {
        bit Z; // Zero
        bit C; // Carry
        bit N; // Negative
        bit V; // Overflow
    } Flags;

endpackage
